module APB_Keyboard(input wire clk,rst_n,
                    input wire );

endmodule